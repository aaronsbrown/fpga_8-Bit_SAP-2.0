import arch_defs_pkg::*;

module control_unit (
    input   wire                                clk,
    input   wire                                reset,
    input   opcode_t                            opcode,
    input   logic           [2:0]               flags,
    output  control_word_t                      control_word
);

    fsm_state_t current_state = S_RESET; // Current microstep in execution
    fsm_state_t next_state = S_RESET; // Next microstep to transition to

    microstep_t current_step; // Current microstep in execution
    microstep_t next_step; // Next microstep to transition to

    logic [1:0] current_byte_count;
    logic [1:0] next_byte_count;
    logic [1:0] num_operand_bytes;
    

    // ==================================================================================================
    // ======================================== ISA OPCODE <=> NUM OPERANDS =============================
    always_comb begin
        num_operand_bytes = 2'bxx;
        case (opcode)
            NOP, HLT: begin
                num_operand_bytes = 2'b00; // No operands
            end
            LDI_A: begin
                num_operand_bytes = 2'b01; // One operand
            end
            LDA: begin
                num_operand_bytes = 2'b10; // One operand
            end
            default: begin
                num_operand_bytes = 2'bxx; // Unknown opcode
                $display($time, " Warning: Unrecognized Opcode %h in case statement", opcode);
            end
        endcase
    end
    
    
    // ==================================================================================================
    // ======================================== SEQ STATE MANAGEMENT =============================
    // Sequential logic for controlling the CPU's operation based on clock and reset signals
    always_ff @(posedge clk) begin 
        if (reset) begin 
            current_state <= S_RESET;
            current_step <= MS0; 
            current_byte_count <= 2'b00; 
        end else begin 
            current_state <= next_state; 
            current_step <= next_step; 
            current_byte_count <= next_byte_count; 
        end
    end

    // ==================================================================================================
    // ======================================== STATE DEFINITION =============================
    // Combinational logic to determine the next state and control word based on the current step
    
    logic check_jump_condition = 1'b0; // Initialize jump condition check
    logic jump_condition_satisfied = 1'b0; // Initialize jump condition satisfied flag
    always_comb begin 

        next_state = current_state;
        next_step = current_step; 
        next_byte_count = current_byte_count;
        control_word = '{default: 0}; 

        case (current_state)
            
            S_RESET: begin
                next_state = S_FETCH_BYTES_0; 
            end
            
            S_FETCH_BYTES_0: begin
                control_word.load_mar_pc = 1'b1; // Load MAR with PC
                next_state = S_FETCH_BYTES_1; 
            end 

            S_FETCH_BYTES_1: begin
                control_word = '{default: 0, oe_ram: 1};
                next_state = S_FETCH_BYTES_2; // Read from RAM
            end

            S_FETCH_BYTES_2: begin
                control_word = '{default: 0, oe_ram: 1, pc_enable: 1};

                if (current_byte_count == 2'b00) begin // opcode
                   control_word.load_ir = 1'b1; // Load instruction register
                end else if ( current_byte_count == 2'b01 ) begin
                    control_word.load_temp_1 = 1'b1; 
                end else if ( current_byte_count == 2'b10 ) begin
                    control_word.load_temp_2 = 1'b1;
                end
                
                next_state = S_WAIT; 
                next_byte_count = current_byte_count + 1; 
            end
            
            S_WAIT: begin
                if ( current_byte_count > num_operand_bytes ) begin
                    next_state = S_EXECUTE;
                    next_byte_count = 2'b00;
                end else begin
                    next_state = S_FETCH_BYTES_0;
                end 
            end
            
            S_EXECUTE: begin
                control_word = microcode_rom[opcode][current_step]; // Fetch control word from microcode ROM
                
                check_jump_condition = control_word.check_zero || control_word.check_carry || control_word.check_negative;
                jump_condition_satisfied = (control_word.check_zero && flags[0]) ||
                                                (control_word.check_carry && flags[1]) ||
                                                (control_word.check_negative && flags[2]);

                if (control_word.halt) begin
                    next_state = S_HALT; 
                    next_step = MS0; 
                // end else if ( check_jump_condition && !jump_condition_satisfied) begin
                   
                //    // Don't Jump! Suppress loading PC with new JMP address if conditions aren't met
                //    control_word.load_pc = 1'b0;
                //    next_state = S_FETCH_0;
                //    next_step = MS0; 
                
                end else if (control_word.last_step) begin
                    next_state = S_FETCH_BYTES_0; 
                    next_step = MS0; 
                end else begin
                    next_state = S_EXECUTE;
                    next_step = current_step + 1; // Increment microstep
                end
            end
            
            S_HALT: begin
                control_word = '{default: 0}; // Default control word
                next_state = S_HALT; // Remain in halt state
            end

            default: begin
                control_word = '{default: 0}; // Default control word
                next_state = S_HALT; // Transition to halt state on error
            end
        endcase
    end

    // ==================================================================================================
    // ======================================== MICROCODE ROM ===========================================
    control_word_t microcode_rom [256][8];
    initial begin
        for (int i = 0; i < 256; i++) begin
            for (int s = 0; s < 8; s++) begin
                microcode_rom[i][s] = '{default: 0}; // Initialize each microstep to zero
            end
        end
        
        // x00
        microcode_rom[NOP][MS0] = '{default: 0, last_step: 1}; 

        // x01
        microcode_rom[HLT][MS0] = '{default: 0, halt: 1}; 

        // x0C
        microcode_rom[LDI_A][MS0] = '{default: 0, oe_temp_1: 1}; 
        microcode_rom[LDI_A][MS1] = '{default: 0, oe_temp_1: 1, load_a: 1, load_flags: 1, last_step: 1}; // todo load_flags, load_sets_zn

    end

endmodule