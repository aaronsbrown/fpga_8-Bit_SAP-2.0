import arch_defs_pkg::*;

module computer (

    input wire clk,
    input wire reset,
    output wire [DATA_WIDTH-1:0] register_OUT,
    output wire cpu_flag_zero_o,
    output wire cpu_flag_carry_o,
    output wire cpu_flag_negative_o,
    output wire [DATA_WIDTH-1:0] cpu_debug_out_B,
    output wire [DATA_WIDTH-1:0] cpu_debug_out_IR,
    output wire [ADDR_WIDTH-1:0] cpu_debug_out_PC
);

    
    logic [ADDR_WIDTH-1:0]  cpu_mem_address;
    logic [DATA_WIDTH-1:0]  cpu_mem_data_out;
    logic [DATA_WIDTH-1:0]  ram_data_out;
    logic                   cpu_mem_write;
    logic                   cpu_mem_read;
    logic                   cpu_load_o;
    logic                   cpu_oe_ram;
    logic                   cpu_oe_a;
    logic [DATA_WIDTH-1:0]  cpu_a_out_bus;
    logic                   cpu_halt;

    cpu u_cpu (
        .clk(clk),
        .reset(reset),
        
        // MEMORY INTERFACE
        .mem_address(cpu_mem_address),
        .mem_read(cpu_mem_read),
        .mem_data_in(ram_data_out),
        .mem_write(cpu_mem_write),
        .mem_data_out(cpu_mem_data_out),
        
        // OUTPUT INTERFACE 
        .load_o(cpu_load_o),
        .oe_ram(cpu_oe_ram),
        .oe_a(cpu_oe_a),
        .a_out_bus(cpu_a_out_bus),

        .halt(cpu_halt),

        // DEBUG SIGNALS
        .flag_zero_o(cpu_flag_zero_o),
        .flag_carry_o(cpu_flag_carry_o),
        .flag_negative_o(cpu_flag_negative_o),
        .debug_out_B(cpu_debug_out_B),
        .debug_out_IR(cpu_debug_out_IR),
        .debug_out_PC(cpu_debug_out_PC)
    );

    ram u_ram (
        .clk(clk),
        .we(cpu_mem_write),
        .address(cpu_mem_address),  
        .data_in(cpu_mem_data_out),
        .data_out(ram_data_out)
    );

    logic [DATA_WIDTH-1:0] register_OUT_data_source;

    assign register_OUT_data_source = 
        (cpu_oe_a) ? cpu_a_out_bus : 
        (cpu_oe_ram) ? ram_data_out : 
        { DATA_WIDTH{1'b0} };


    register_nbit #( .N(DATA_WIDTH) ) u_register_OUT (
        .clk(clk),
        .reset(reset),
        .load(cpu_load_o),
        .data_in(register_OUT_data_source),
        .latched_data(register_OUT)
    );

endmodule